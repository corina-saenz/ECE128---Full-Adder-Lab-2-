`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/09/2025 02:07:15 PM
// Design Name: 
// Module Name: tb_fa1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_fa1(
    input [3:0] swA,
    input [3:0] swB,
    input swCI,
    input [3:0] ledSUM,
    input ledCO
    );
endmodule
